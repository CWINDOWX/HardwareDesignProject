`timescale 1ns / 1ps

/*
 * Branch_Cmp.v
 * ��֧�Ƚ��� - �Ƚ������Ĵ�����ֵ���жϷ�֧�Ƿ����
 * Member 4: ��Ա4
 */

module Branch_Cmp(
    input  [31:0] a,          // ��һ����������rs��
    input  [31:0] b,          // �ڶ�����������rt��
    input  [2:0]  cmp_op,     // �Ƚϲ�������
    output reg    cmp_result  // �ȽϽ����1:��֧, 0:����֧��
);

// �Ƚϲ������壺
// 000: BEQ  - ������֧ (a == b)
// 001: BNE  - �������֧ (a != b)
// 010: BGTZ - ����0���֧ (a > 0)
// 011: BLEZ - С�ڵ���0���֧ (a <= 0)
// 100: BLTZ - С��0���֧ (a < 0)
// 101: BGEZ - ���ڵ���0���֧ (a >= 0)

always @(*) begin
    case (cmp_op)
        3'b000:  cmp_result = (a == b);                           // BEQ
        3'b001:  cmp_result = (a != b);                           // BNE
        3'b010:  cmp_result = (~a[31]) & (a != 32'h00000000);    // BGTZ: �����ҷ�0
        3'b011:  cmp_result = a[31] | (a == 32'h00000000);       // BLEZ: ������0
        3'b100:  cmp_result = a[31];                             // BLTZ: ����λ=1
        3'b101:  cmp_result = ~a[31];                            // BGEZ: ����λ=0
        default: cmp_result = 1'b0;
    endcase
end

endmodule